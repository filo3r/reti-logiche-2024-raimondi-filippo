-------------------------------------------------------------------------
-- Prova Finale di Reti Logiche                                        --
-- Anno Accademico 2023-2024                                           --
-- Politecnico di Milano                                               --
-- Filippo Raimondi                                                    --
-- 10809051                                                            --
-- Testbench 4: K = 1023                                               --
-------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;

ENTITY project_tb_4 IS
END project_tb_4;

ARCHITECTURE project_tb_4_arch OF project_tb_4 IS

    -- Costanti
    CONSTANT CLOCK_PERIOD : TIME := 20 ns;
    CONSTANT SCENARIO_ADDRESS : INTEGER := 40000;
    CONSTANT SCENARIO_LENGTH : INTEGER := 1023;

    -- Tipi custom
    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    TYPE scenario_type IS ARRAY (0 TO SCENARIO_LENGTH * 2 - 1) OF INTEGER;

    -- Segnali principali
    SIGNAL tb_clk         : STD_LOGIC := '0';
    SIGNAL tb_rst         : STD_LOGIC;
    SIGNAL tb_start       : STD_LOGIC;
    SIGNAL tb_done        : STD_LOGIC;
    SIGNAL tb_add         : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL tb_k           : STD_LOGIC_VECTOR(9 DOWNTO 0);

    SIGNAL tb_o_mem_addr  : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL tb_o_mem_data  : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL tb_i_mem_data  : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL tb_o_mem_we    : STD_LOGIC;
    SIGNAL tb_o_mem_en    : STD_LOGIC;

    SIGNAL exc_o_mem_addr : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL exc_o_mem_data : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL exc_o_mem_we   : STD_LOGIC;
    SIGNAL exc_o_mem_en   : STD_LOGIC;

    SIGNAL init_o_mem_addr : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL init_o_mem_data : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL init_o_mem_we   : STD_LOGIC;
    SIGNAL init_o_mem_en   : STD_LOGIC;

    SIGNAL memory_control : STD_LOGIC := '0';
    SIGNAL RAM            : ram_type := (OTHERS => "00000000");

    SIGNAL scenario_input : scenario_type := (86, 0, 0, 0, 0, 0, 0, 0, 74, 0, 0, 0, 42, 0, 0, 0, 121, 0, 58, 0, 0, 0, 0, 0, 127, 0, 199, 0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
                                              239, 0, 224, 0, 0, 0, 0, 0, 227, 0, 0, 0, 0, 0, 83, 0, 78, 0, 0, 0, 150, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 0, 25, 0, 213, 0, 19, 0, 
                                              72, 0, 196, 0, 213, 0, 0, 0, 0, 0, 231, 0, 21, 0, 0, 0, 196, 0, 0, 0, 165, 0, 0, 0, 0, 0, 89, 0, 0, 0, 15, 0, 0, 0, 123, 0, 0, 0, 
                                              89, 0, 0, 0, 179, 0, 191, 0, 120, 0, 0, 0, 0, 0, 74, 0, 24, 0, 0, 0, 40, 0, 0, 0, 0, 0, 132, 0, 0, 0, 180, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
                                              235, 0, 0, 0, 14, 0, 92, 0, 0, 0, 0, 0, 116, 0, 51, 0, 0, 0, 0, 0, 196, 0, 123, 0, 239, 0, 227, 0, 0, 0, 244, 0, 74, 0, 0, 0, 0, 0, 0, 0, 
                                              177, 0, 0, 0, 100, 0, 28, 0, 0, 0, 0, 0, 0, 0, 131, 0, 0, 0, 0, 0, 0, 0, 0, 0, 248, 0, 152, 0, 231, 0, 0, 0, 19, 0, 225, 0, 159, 0, 0, 0, 
                                              0, 0, 0, 0, 0, 0, 176, 0, 196, 0, 71, 0, 0, 0, 1, 0, 9, 0, 0, 0, 0, 0, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 201, 0, 41, 0, 0, 0, 114, 0, 0, 
                                              0, 0, 0, 181, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 211, 0, 0, 0, 138, 0, 0, 0, 32, 0, 0, 0, 90, 0, 137, 0, 176, 0, 0, 0, 
                                              218, 0, 0, 0, 145, 0, 5, 0, 0, 0, 0, 0, 128, 0, 37, 0, 0, 0, 12, 0, 159, 0, 0, 0, 210, 0, 231, 0, 160, 0, 0, 0, 177, 0, 112, 0, 188, 0, 37, 0, 
                                              0, 0, 226, 0, 0, 0, 9, 0, 143, 0, 0, 0, 224, 0, 221, 0, 0, 0, 205, 0, 0, 0, 0, 0, 199, 0, 250, 0, 6, 0, 130, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
                                              0, 230, 0, 0, 0, 0, 0, 0, 0, 253, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 187, 0, 63, 0, 174, 0, 114, 0, 0, 0, 103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
                                              84, 0, 58, 0, 0, 0, 155, 0, 0, 0, 133, 0, 27, 0, 4, 0, 32, 0, 151, 0, 148, 0, 175, 0, 0, 0, 0, 0, 52, 0, 64, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
                                              124, 0, 243, 0, 111, 0, 0, 0, 220, 0, 39, 0, 177, 0, 0, 0, 9, 0, 11, 0, 0, 0, 180, 0, 184, 0, 94, 0, 0, 0, 203, 0, 0, 0, 173, 0, 0, 0, 108, 0, 
                                              169, 0, 0, 0, 137, 0, 30, 0, 0, 0, 202, 0, 63, 0, 0, 0, 78, 0, 159, 0, 0, 0, 36, 0, 0, 0, 78, 0, 248, 0, 0, 0, 0, 0, 39, 0, 94, 0, 195, 0, 0, 0, 
                                              101, 0, 0, 0, 91, 0, 0, 0, 221, 0, 2, 0, 215, 0, 0, 0, 240, 0, 40, 0, 0, 0, 180, 0, 0, 0, 152, 0, 0, 0, 0, 0, 3, 0, 197, 0, 0, 0, 165, 0, 0, 0, 0, 
                                              0, 195, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 251, 0, 89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 221, 0, 0, 0, 0, 0, 0, 0, 245, 0, 0, 0, 75, 0, 0, 0, 
                                              0, 0, 0, 0, 0, 0, 92, 0, 0, 0, 0, 0, 175, 0, 117, 0, 104, 0, 129, 0, 0, 0, 0, 0, 148, 0, 212, 0, 159, 0, 135, 0, 0, 0, 174, 0, 0, 0, 16, 0, 128, 
                                              0, 42, 0, 0, 0, 220, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 253, 0, 4, 0, 0, 0, 24, 0, 0, 0, 0, 0, 99, 0, 0, 0, 232, 0, 
                                              66, 0, 0, 0, 0, 0, 196, 0, 0, 0, 0, 0, 238, 0, 30, 0, 14, 0, 0, 0, 0, 0, 0, 0, 92, 0, 98, 0, 95, 0, 193, 0, 65, 0, 0, 0, 87, 0, 247, 0, 0, 0, 0, 
                                              0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 62, 0, 177, 0, 0, 0, 0, 0, 0, 0, 92, 0, 0, 0, 204, 0, 28, 0, 0, 0, 53, 0, 0, 0, 250, 0, 
                                              0, 0, 64, 0, 6, 0, 208, 0, 60, 0, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 221, 0, 205, 0, 83, 0, 0, 0, 0, 0, 115, 0, 0, 0, 113, 0, 0, 0, 25, 0, 162, 0, 0, 
                                              0, 189, 0, 0, 0, 0, 0, 167, 0, 190, 0, 0, 0, 0, 0, 0, 0, 5, 0, 43, 0, 106, 0, 0, 0, 171, 0, 0, 0, 33, 0, 94, 0, 0, 0, 0, 0, 162, 0, 133, 0, 134, 
                                              0, 118, 0, 215, 0, 0, 0, 127, 0, 113, 0, 0, 0, 79, 0, 116, 0, 0, 0, 20, 0, 0, 0, 6, 0, 0, 0, 235, 0, 127, 0, 7, 0, 129, 0, 0, 0, 0, 0, 0, 0, 0, 0,
                                              0, 0, 238, 0, 253, 0, 140, 0, 0, 0, 0, 0, 90, 0, 0, 0, 0, 0, 0, 0, 207, 0, 0, 0, 0, 0, 0, 0, 202, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 253, 0, 0, 0, 
                                              185, 0, 0, 0, 0, 0, 0, 0, 247, 0, 0, 0, 0, 0, 0, 0, 0, 0, 255, 0, 223, 0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 152, 0, 0, 0, 162, 0, 6, 0, 50, 
                                              0, 148, 0, 0, 0, 92, 0, 219, 0, 90, 0, 0, 0, 0, 0, 205, 0, 0, 0, 0, 0, 142, 0, 0, 0, 0, 0, 209, 0, 0, 0, 148, 0, 249, 0, 22, 0, 0, 0, 90, 0, 0, 0, 0, 
                                              0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112, 0, 0, 0, 44, 0, 76, 0, 31, 0, 0, 0, 0, 0, 151, 0, 0, 0, 148, 0, 45, 0, 99, 0, 43, 0, 198, 0, 
                                              0, 0, 129, 0, 53, 0, 0, 0, 172, 0, 186, 0, 46, 0, 209, 0, 0, 0, 124, 0, 87, 0, 0, 0, 0, 0, 175, 0, 22, 0, 26, 0, 157, 0, 0, 0, 170, 0, 0, 0, 0, 0, 28, 
                                              0, 230, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 12, 0, 68, 0, 0, 0, 41, 0, 244, 0, 24, 0, 0, 0, 0, 0, 38, 0, 1, 0, 160, 0, 62, 0, 33, 0, 0, 0, 61, 0, 44, 0, 
                                              34, 0, 194, 0, 66, 0, 141, 0, 0, 0, 85, 0, 0, 0, 104, 0, 0, 0, 68, 0, 0, 0, 60, 0, 0, 0, 119, 0, 42, 0, 214, 0, 0, 0, 50, 0, 0, 0, 167, 0, 87, 0, 0, 0, 
                                              0, 0, 88, 0, 103, 0, 227, 0, 121, 0, 0, 0, 28, 0, 28, 0, 0, 0, 163, 0, 0, 0, 180, 0, 215, 0, 49, 0, 33, 0, 176, 0, 22, 0, 0, 0, 14, 0, 192, 0, 97, 0, 0, 0, 
                                              173, 0, 234, 0, 94, 0, 0, 0, 0, 0, 0, 0, 56, 0, 139, 0, 133, 0, 0, 0, 61, 0, 0, 0, 124, 0, 34, 0, 116, 0, 0, 0, 0, 0, 44, 0, 0, 0, 169, 0, 0, 0, 0, 0, 
                                              211, 0, 129, 0, 0, 0, 0, 0, 135, 0, 0, 0, 167, 0, 133, 0, 0, 0, 64, 0, 0, 0, 34, 0, 0, 0, 2, 0, 0, 0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 0, 0, 0, 214, 0, 
                                              76, 0, 0, 0, 0, 0, 132, 0, 103, 0, 66, 0, 207, 0, 0, 0, 0, 0, 0, 0, 0, 0, 217, 0, 30, 0, 166, 0, 217, 0, 220, 0, 31, 0, 0, 0, 0, 0, 85, 0, 0, 0, 0, 0, 
                                              0, 0, 250, 0, 0, 0, 147, 0, 0, 0, 88, 0, 77, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 249, 0, 0, 0, 0, 0, 0, 0, 151, 0, 169, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
                                              0, 0, 242, 0, 254, 0, 0, 0, 0, 0, 245, 0, 0, 0, 0, 0, 0, 0, 142, 0, 0, 0, 15, 0, 0, 0, 0, 0, 207, 0, 248, 0, 0, 0, 163, 0, 0, 0, 232, 0, 60, 0, 98, 0, 
                                              0, 0, 0, 0, 41, 0, 8, 0, 196, 0, 0, 0, 195, 0, 0, 0, 0, 0, 73, 0, 0, 0, 0, 0, 202, 0, 169, 0, 86, 0, 0, 0, 233, 0, 0, 0, 92, 0, 51, 0, 0, 0, 0, 0, 91, 
                                              0, 44, 0, 0, 0, 0, 0, 0, 0, 52, 0, 0, 0, 135, 0, 76, 0, 0, 0, 176, 0, 0, 0, 0, 0, 57, 0, 0, 0, 84, 0, 0, 0, 250, 0, 0, 0, 100, 0, 0, 0, 0, 0, 0, 0, 0, 
                                              0, 0, 0, 93, 0, 71, 0, 0, 0, 134, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 136, 0, 0, 0, 0, 0, 22, 0, 53, 0, 0, 0, 0, 
                                              0, 186, 0, 245, 0, 189, 0, 217, 0, 0, 0, 0, 0, 100, 0, 0, 0, 0, 0, 178, 0, 0, 0, 188, 0, 0, 0, 0, 0, 0, 0, 191, 0, 4, 0, 42, 0, 0, 0, 117, 0, 0, 0, 0, 0, 
                                              0, 0, 0, 0, 148, 0, 101, 0, 0, 0, 87, 0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 50, 0, 102, 0, 255, 0, 0, 
                                              0, 0, 0, 0, 0, 109, 0, 0, 0, 47, 0, 0, 0, 151, 0, 241, 0, 0, 0, 0, 0, 0, 0, 141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 66, 0, 0, 0, 81, 0, 247, 0, 0, 0, 239, 
                                              0, 0, 0, 128, 0, 55, 0, 209, 0, 0, 0, 108, 0, 0, 0, 0, 0, 205, 0, 56, 0, 210, 0, 0, 0, 122, 0, 1, 0, 0, 0, 72, 0, 86, 0, 128, 0, 60, 0, 4, 0, 44, 0, 0, 0, 
                                              110, 0, 88, 0, 0, 0, 0, 0, 46, 0, 82, 0, 0, 0, 9, 0, 209, 0, 175, 0, 0, 0, 155, 0, 171, 0, 0, 0, 0, 0, 0, 0, 182, 0, 32, 0, 162, 0, 9, 0, 0, 0, 255, 0, 64, 
                                              0, 0, 0, 0, 0, 21, 0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 172, 0, 0, 0, 201, 0, 0, 0, 0, 0, 0, 0, 185, 0, 89, 0, 0, 0, 0, 0, 117, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
                                              73, 0, 0, 0, 142, 0, 23, 0, 99, 0, 240, 0, 214, 0, 232, 0, 171, 0, 12, 0, 172, 0, 204, 0, 216, 0, 148, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 0, 234, 0, 0, 0, 0, 0, 
                                              73, 0, 0, 0, 0, 0, 50, 0, 0, 0, 214, 0, 0, 0, 0, 0, 138, 0, 0, 0, 184, 0, 0, 0, 31, 0, 0, 0, 0, 0, 71, 0, 0, 0, 0, 0, 164, 0, 127, 0, 0, 0, 0, 0, 169, 0);

    SIGNAL scenario_full : scenario_type := (86, 31, 86, 30, 86, 29, 86, 28, 74, 31, 74, 30, 42, 31, 42, 30, 121, 31, 58, 31, 58, 30, 58, 29, 127, 31, 199, 31, 199, 30, 55, 31, 55, 30, 55, 29, 
                                             55, 28, 55, 27, 239, 31, 224, 31, 224, 30, 224, 29, 227, 31, 227, 30, 227, 29, 83, 31, 78, 31, 78, 30, 150, 31, 150, 30, 150, 29, 150, 28, 150, 27, 
                                             67, 31, 25, 31, 213, 31, 19, 31, 72, 31, 196, 31, 213, 31, 213, 30, 213, 29, 231, 31, 21, 31, 21, 30, 196, 31, 196, 30, 165, 31, 165, 30, 165, 29, 89, 
                                             31, 89, 30, 15, 31, 15, 30, 123, 31, 123, 30, 89, 31, 89, 30, 179, 31, 191, 31, 120, 31, 120, 30, 120, 29, 74, 31, 24, 31, 24, 30, 40, 31, 40, 30, 40, 
                                             29, 132, 31, 132, 30, 180, 31, 180, 30, 180, 29, 180, 28, 180, 27, 235, 31, 235, 30, 14, 31, 92, 31, 92, 30, 92, 29, 116, 31, 51, 31, 51, 30, 51, 29, 
                                             196, 31, 123, 31, 239, 31, 227, 31, 227, 30, 244, 31, 74, 31, 74, 30, 74, 29, 74, 28, 177, 31, 177, 30, 100, 31, 28, 31, 28, 30, 28, 29, 28, 28, 131, 
                                             31, 131, 30, 131, 29, 131, 28, 131, 27, 248, 31, 152, 31, 231, 31, 231, 30, 19, 31, 225, 31, 159, 31, 159, 30, 159, 29, 159, 28, 159, 27, 176, 31, 
                                             196, 31, 71, 31, 71, 30, 1, 31, 9, 31, 9, 30, 9, 29, 81, 31, 81, 30, 81, 29, 81, 28, 81, 27, 81, 26, 201, 31, 41, 31, 41, 30, 114, 31, 114, 30, 114, 29, 
                                             181, 31, 181, 30, 181, 29, 181, 28, 181, 27, 181, 26, 181, 25, 181, 24, 181, 23, 181, 22, 211, 31, 211, 30, 138, 31, 138, 30, 32, 31, 32, 30, 90, 31, 137, 
                                             31, 176, 31, 176, 30, 218, 31, 218, 30, 145, 31, 5, 31, 5, 30, 5, 29, 128, 31, 37, 31, 37, 30, 12, 31, 159, 31, 159, 30, 210, 31, 231, 31, 160, 31, 160, 30, 
                                             177, 31, 112, 31, 188, 31, 37, 31, 37, 30, 226, 31, 226, 30, 9, 31, 143, 31, 143, 30, 224, 31, 221, 31, 221, 30, 205, 31, 205, 30, 205, 29, 199, 31, 250, 31, 
                                             6, 31, 130, 31, 130, 30, 130, 29, 130, 28, 130, 27, 130, 26, 130, 25, 230, 31, 230, 30, 230, 29, 230, 28, 253, 31, 43, 31, 43, 30, 43, 29, 43, 28, 43, 27, 187, 
                                             31, 63, 31, 174, 31, 114, 31, 114, 30, 103, 31, 103, 30, 103, 29, 103, 28, 103, 27, 103, 26, 84, 31, 58, 31, 58, 30, 155, 31, 155, 30, 133, 31, 27, 31, 4, 31, 
                                             32, 31, 151, 31, 148, 31, 175, 31, 175, 30, 175, 29, 52, 31, 64, 31, 43, 31, 43, 30, 43, 29, 43, 28, 43, 27, 124, 31, 243, 31, 111, 31, 111, 30, 220, 31, 39, 31, 
                                             177, 31, 177, 30, 9, 31, 11, 31, 11, 30, 180, 31, 184, 31, 94, 31, 94, 30, 203, 31, 203, 30, 173, 31, 173, 30, 108, 31, 169, 31, 169, 30, 137, 31, 30, 31, 30, 
                                             30, 202, 31, 63, 31, 63, 30, 78, 31, 159, 31, 159, 30, 36, 31, 36, 30, 78, 31, 248, 31, 248, 30, 248, 29, 39, 31, 94, 31, 195, 31, 195, 30, 101, 31, 101, 30, 
                                             91, 31, 91, 30, 221, 31, 2, 31, 215, 31, 215, 30, 240, 31, 40, 31, 40, 30, 180, 31, 180, 30, 152, 31, 152, 30, 152, 29, 3, 31, 197, 31, 197, 30, 165, 31, 165, 
                                             30, 165, 29, 195, 31, 195, 30, 195, 29, 195, 28, 195, 27, 195, 26, 251, 31, 89, 31, 89, 30, 89, 29, 89, 28, 89, 27, 89, 26, 89, 25, 221, 31, 221, 30, 221, 29, 
                                             221, 28, 245, 31, 245, 30, 75, 31, 75, 30, 75, 29, 75, 28, 75, 27, 92, 31, 92, 30, 92, 29, 175, 31, 117, 31, 104, 31, 129, 31, 129, 30, 129, 29, 148, 31, 212, 
                                             31, 159, 31, 135, 31, 135, 30, 174, 31, 174, 30, 16, 31, 128, 31, 42, 31, 42, 30, 220, 31, 220, 30, 220, 29, 220, 28, 220, 27, 220, 26, 220, 25, 220, 24, 220, 
                                             23, 220, 22, 220, 21, 253, 31, 4, 31, 4, 30, 24, 31, 24, 30, 24, 29, 99, 31, 99, 30, 232, 31, 66, 31, 66, 30, 66, 29, 196, 31, 196, 30, 196, 29, 238, 31, 30, 
                                             31, 14, 31, 14, 30, 14, 29, 14, 28, 92, 31, 98, 31, 95, 31, 193, 31, 65, 31, 65, 30, 87, 31, 247, 31, 247, 30, 247, 29, 247, 28, 247, 27, 247, 26, 247, 25, 
                                             247, 24, 247, 23, 247, 22, 19, 31, 19, 30, 62, 31, 177, 31, 177, 30, 177, 29, 177, 28, 92, 31, 92, 30, 204, 31, 28, 31, 28, 30, 53, 31, 53, 30, 250, 31, 
                                             250, 30, 64, 31, 6, 31, 208, 31, 60, 31, 76, 31, 76, 30, 76, 29, 76, 28, 76, 27, 221, 31, 205, 31, 83, 31, 83, 30, 83, 29, 115, 31, 115, 30, 113, 31, 113, 
                                             30, 25, 31, 162, 31, 162, 30, 189, 31, 189, 30, 189, 29, 167, 31, 190, 31, 190, 30, 190, 29, 190, 28, 5, 31, 43, 31, 106, 31, 106, 30, 171, 31, 171, 30, 33, 
                                             31, 94, 31, 94, 30, 94, 29, 162, 31, 133, 31, 134, 31, 118, 31, 215, 31, 215, 30, 127, 31, 113, 31, 113, 30, 79, 31, 116, 31, 116, 30, 20, 31, 20, 30, 6, 31, 
                                             6, 30, 235, 31, 127, 31, 7, 31, 129, 31, 129, 30, 129, 29, 129, 28, 129, 27, 129, 26, 238, 31, 253, 31, 140, 31, 140, 30, 140, 29, 90, 31, 90, 30, 90, 29, 90, 
                                             28, 207, 31, 207, 30, 207, 29, 207, 28, 202, 31, 35, 31, 35, 30, 35, 29, 35, 28, 35, 27, 253, 31, 253, 30, 185, 31, 185, 30, 185, 29, 185, 28, 247, 31, 247, 
                                             30, 247, 29, 247, 28, 247, 27, 255, 31, 223, 31, 223, 30, 55, 31, 55, 30, 55, 29, 55, 28, 22, 31, 22, 30, 152, 31, 152, 30, 162, 31, 6, 31, 50, 31, 148, 31, 
                                             148, 30, 92, 31, 219, 31, 90, 31, 90, 30, 90, 29, 205, 31, 205, 30, 205, 29, 142, 31, 142, 30, 142, 29, 209, 31, 209, 30, 148, 31, 249, 31, 22, 31, 22, 30, 
                                             90, 31, 90, 30, 90, 29, 90, 28, 90, 27, 90, 26, 90, 25, 90, 24, 90, 23, 90, 22, 90, 21, 112, 31, 112, 30, 44, 31, 76, 31, 31, 31, 31, 30, 31, 29, 151, 31, 
                                             151, 30, 148, 31, 45, 31, 99, 31, 43, 31, 198, 31, 198, 30, 129, 31, 53, 31, 53, 30, 172, 31, 186, 31, 46, 31, 209, 31, 209, 30, 124, 31, 87, 31, 87, 30, 
                                             87, 29, 175, 31, 22, 31, 26, 31, 157, 31, 157, 30, 170, 31, 170, 30, 170, 29, 28, 31, 230, 31, 230, 30, 230, 29, 230, 28, 30, 31, 30, 30, 12, 31, 68, 31, 
                                             68, 30, 41, 31, 244, 31, 24, 31, 24, 30, 24, 29, 38, 31, 1, 31, 160, 31, 62, 31, 33, 31, 33, 30, 61, 31, 44, 31, 34, 31, 194, 31, 66, 31, 141, 31, 141, 
                                             30, 85, 31, 85, 30, 104, 31, 104, 30, 68, 31, 68, 30, 60, 31, 60, 30, 119, 31, 42, 31, 214, 31, 214, 30, 50, 31, 50, 30, 167, 31, 87, 31, 87, 30, 87, 29, 
                                             88, 31, 103, 31, 227, 31, 121, 31, 121, 30, 28, 31, 28, 31, 28, 30, 163, 31, 163, 30, 180, 31, 215, 31, 49, 31, 33, 31, 176, 31, 22, 31, 22, 30, 14, 31, 
                                             192, 31, 97, 31, 97, 30, 173, 31, 234, 31, 94, 31, 94, 30, 94, 29, 94, 28, 56, 31, 139, 31, 133, 31, 133, 30, 61, 31, 61, 30, 124, 31, 34, 31, 116, 31, 
                                             116, 30, 116, 29, 44, 31, 44, 30, 169, 31, 169, 30, 169, 29, 211, 31, 129, 31, 129, 30, 129, 29, 135, 31, 135, 30, 167, 31, 133, 31, 133, 30, 64, 31, 
                                             64, 30, 34, 31, 34, 30, 2, 31, 2, 30, 63, 31, 63, 30, 63, 29, 63, 28, 63, 27, 54, 31, 54, 30, 214, 31, 76, 31, 76, 30, 76, 29, 132, 31, 103, 31, 66, 
                                             31, 207, 31, 207, 30, 207, 29, 207, 28, 207, 27, 217, 31, 30, 31, 166, 31, 217, 31, 220, 31, 31, 31, 31, 30, 31, 29, 85, 31, 85, 30, 85, 29, 85, 28, 
                                             250, 31, 250, 30, 147, 31, 147, 30, 88, 31, 77, 31, 43, 31, 43, 30, 43, 29, 43, 28, 43, 27, 249, 31, 249, 30, 249, 29, 249, 28, 151, 31, 169, 31, 169, 
                                             30, 169, 29, 169, 28, 169, 27, 169, 26, 169, 25, 242, 31, 254, 31, 254, 30, 254, 29, 245, 31, 245, 30, 245, 29, 245, 28, 142, 31, 142, 30, 15, 31, 15, 
                                             30, 15, 29, 207, 31, 248, 31, 248, 30, 163, 31, 163, 30, 232, 31, 60, 31, 98, 31, 98, 30, 98, 29, 41, 31, 8, 31, 196, 31, 196, 30, 195, 31, 195, 30, 
                                             195, 29, 73, 31, 73, 30, 73, 29, 202, 31, 169, 31, 86, 31, 86, 30, 233, 31, 233, 30, 92, 31, 51, 31, 51, 30, 51, 29, 91, 31, 44, 31, 44, 30, 44, 29, 
                                             44, 28, 52, 31, 52, 30, 135, 31, 76, 31, 76, 30, 176, 31, 176, 30, 176, 29, 57, 31, 57, 30, 84, 31, 84, 30, 250, 31, 250, 30, 100, 31, 100, 30, 100, 
                                             29, 100, 28, 100, 27, 100, 26, 93, 31, 71, 31, 71, 30, 134, 31, 15, 31, 15, 30, 15, 29, 15, 28, 15, 27, 15, 26, 33, 31, 33, 30, 33, 29, 33, 28, 33, 
                                             27, 33, 26, 136, 31, 136, 30, 136, 29, 22, 31, 53, 31, 53, 30, 53, 29, 186, 31, 245, 31, 189, 31, 217, 31, 217, 30, 217, 29, 100, 31, 100, 30, 100, 
                                             29, 178, 31, 178, 30, 188, 31, 188, 30, 188, 29, 188, 28, 191, 31, 4, 31, 42, 31, 42, 30, 117, 31, 117, 30, 117, 29, 117, 28, 117, 27, 148, 31, 101, 
                                             31, 101, 30, 87, 31, 87, 30, 37, 31, 37, 30, 37, 29, 37, 28, 149, 31, 149, 30, 149, 29, 149, 28, 149, 27, 149, 26, 9, 31, 9, 30, 9, 29, 50, 31, 102, 
                                             31, 255, 31, 255, 30, 255, 29, 255, 28, 109, 31, 109, 30, 47, 31, 47, 30, 151, 31, 241, 31, 241, 30, 241, 29, 241, 28, 141, 31, 141, 30, 141, 29, 
                                             141, 28, 141, 27, 31, 31, 66, 31, 66, 30, 81, 31, 247, 31, 247, 30, 239, 31, 239, 30, 128, 31, 55, 31, 209, 31, 209, 30, 108, 31, 108, 30, 108, 
                                             29, 205, 31, 56, 31, 210, 31, 210, 30, 122, 31, 1, 31, 1, 30, 72, 31, 86, 31, 128, 31, 60, 31, 4, 31, 44, 31, 44, 30, 110, 31, 88, 31, 88, 30, 
                                             88, 29, 46, 31, 82, 31, 82, 30, 9, 31, 209, 31, 175, 31, 175, 30, 155, 31, 171, 31, 171, 30, 171, 29, 171, 28, 182, 31, 32, 31, 162, 31, 9, 31, 
                                             9, 30, 255, 31, 64, 31, 64, 30, 64, 29, 21, 31, 21, 30, 37, 31, 37, 30, 37, 29, 37, 28, 37, 27, 172, 31, 172, 30, 201, 31, 201, 30, 201, 29, 201, 
                                             28, 185, 31, 89, 31, 89, 30, 89, 29, 117, 31, 117, 30, 117, 29, 117, 28, 117, 27, 73, 31, 73, 30, 142, 31, 23, 31, 99, 31, 240, 31, 214, 31, 232, 
                                             31, 171, 31, 12, 31, 172, 31, 204, 31, 216, 31, 148, 31, 148, 30, 148, 29, 46, 31, 46, 30, 46, 29, 234, 31, 234, 30, 234, 29, 73, 31, 73, 30, 73, 
                                             29, 50, 31, 50, 30, 214, 31, 214, 30, 214, 29, 138, 31, 138, 30, 184, 31, 184, 30, 31, 31, 31, 30, 31, 29, 71, 31, 71, 30, 71, 29, 164, 31, 127, 31, 
                                             127, 30, 127, 29, 169, 31);

    -- Componenti
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk      : IN  STD_LOGIC;
            i_rst      : IN  STD_LOGIC;
            i_start    : IN  STD_LOGIC;
            i_add      : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_k        : IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
            o_done     : OUT STD_LOGIC;
            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_data : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we   : OUT STD_LOGIC;
            o_mem_en   : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN

    -- Instanza del DUT
    UUT : project_reti_logiche
        PORT MAP (
            i_clk      => tb_clk,
            i_rst      => tb_rst,
            i_start    => tb_start,
            i_add      => tb_add,
            i_k        => tb_k,
            o_done     => tb_done,
            o_mem_addr => exc_o_mem_addr,
            i_mem_data => tb_i_mem_data,
            o_mem_data => exc_o_mem_data,
            o_mem_we   => exc_o_mem_we,
            o_mem_en   => exc_o_mem_en
        );

    -- Generazione del clock
    tb_clk <= NOT tb_clk AFTER CLOCK_PERIOD / 2;

    -- Comportamento della memoria
    MEM : PROCESS(tb_clk)
    BEGIN
        IF tb_clk'EVENT AND tb_clk = '1' THEN
            IF tb_o_mem_en = '1' THEN
                IF tb_o_mem_we = '1' THEN
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data AFTER 1 ns;
                    tb_i_mem_data <= tb_o_mem_data AFTER 1 ns;
                ELSE
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) AFTER 1 ns;
                END IF;
            END IF;
        END IF;
    END PROCESS;

    -- Scambio segnali memoria
    memory_signal_swapper : PROCESS(memory_control, init_o_mem_addr, init_o_mem_data, init_o_mem_en, init_o_mem_we, 
                                    exc_o_mem_addr, exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    BEGIN
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        IF memory_control = '1' THEN
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        END IF;
    END PROCESS;

    -- Generazione scenario iniziale
    create_scenario : PROCESS
    BEGIN
        WAIT FOR 50 ns;

        -- Inizializzazione segnali e reset del componente
        tb_start <= '0';
        tb_add <= (OTHERS => '0');
        tb_k   <= (OTHERS => '0');
        tb_rst <= '1';

        -- Attendere un po' di tempo per il reset
        WAIT FOR 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memoria controllata dal testbench

        -- Skew dei segnali del testbench rispetto al clock
        WAIT UNTIL FALLING_EDGE(tb_clk);

        -- Configurazione della memoria
        FOR i IN 0 TO SCENARIO_LENGTH * 2 - 1 LOOP
            init_o_mem_addr <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS + i, 16));
            init_o_mem_data <= std_logic_vector(to_unsigned(scenario_input(i), 8));
            init_o_mem_en   <= '1';
            init_o_mem_we   <= '1';
            WAIT UNTIL RISING_EDGE(tb_clk);
        END LOOP;

        WAIT UNTIL FALLING_EDGE(tb_clk);

        -- Passaggio del controllo memoria al componente
        memory_control <= '1';

        -- Configurazione dei segnali di input per il componente
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        tb_start <= '1';

        -- Attendere che il componente completi l'elaborazione
        WHILE tb_done /= '1' LOOP
            WAIT UNTIL RISING_EDGE(tb_clk);
        END LOOP;

        -- Disabilitazione di start
        WAIT FOR 5 ns;
        tb_start <= '0';

        WAIT; -- Terminazione della simulazione
    END PROCESS;

        -- Routine di verifica
        test_routine : PROCESS
        BEGIN
            -- Attendere l'attivazione del reset
            WAIT UNTIL tb_rst = '1';
            WAIT FOR 25 ns;
    
            -- Verifica: o_done deve essere '0' durante il reset
            ASSERT tb_done = '0' REPORT "TEST FALLITO: o_done != 0 durante reset" SEVERITY FAILURE;
    
            -- Attendere la disattivazione del reset
            WAIT UNTIL tb_rst = '0';
    
            -- Verifica: o_done deve essere '0' dopo il reset e prima dello start
            WAIT UNTIL FALLING_EDGE(tb_clk);
            ASSERT tb_done = '0' REPORT "TEST FALLITO: o_done != 0 dopo reset prima di start" SEVERITY FAILURE;
    
            -- Attendere l'attivazione del segnale di start
            WAIT UNTIL RISING_EDGE(tb_start);
    
            -- Attendere il completamento del componente
            WHILE tb_done /= '1' LOOP
                WAIT UNTIL RISING_EDGE(tb_clk);
            END LOOP;
    
            -- Verifica: dopo il completamento, la memoria non deve essere scritta
            ASSERT tb_o_mem_en = '0' OR tb_o_mem_we = '0' REPORT "TEST FALLITO: o_mem_en != 0, la memoria non dovrebbe essere scritta dopo il completamento" SEVERITY FAILURE;
    
            -- Verifica: il contenuto della RAM corrisponde ai dati attesi
            FOR i IN 0 TO SCENARIO_LENGTH * 2 - 1 LOOP
                ASSERT RAM(SCENARIO_ADDRESS + i) = std_logic_vector(to_unsigned(scenario_full(i), 8)) REPORT "TEST FALLITO: OFFSET = " & INTEGER'IMAGE(i) & " ATTESO = " & INTEGER'IMAGE(scenario_full(i)) & " TROVATO = " & INTEGER'IMAGE(to_integer(unsigned(RAM(SCENARIO_ADDRESS + i)))) SEVERITY FAILURE;
            END LOOP;
    
            -- Attendere la disattivazione di start
            WAIT UNTIL FALLING_EDGE(tb_start);
    
            -- Verifica: o_done deve rimanere '1' dopo il completamento
            ASSERT tb_done = '1' REPORT "TEST FALLITO: o_done != 0 dopo reset prima di start" SEVERITY FAILURE;
    
            -- Attendere il termine del segnale o_done
            WAIT UNTIL FALLING_EDGE(tb_done);
    
            -- Segnalazione di successo della simulazione
            ASSERT FALSE REPORT "Simulazione completata! TEST PASSATO" SEVERITY FAILURE;
        END PROCESS;
    
END ARCHITECTURE;